library verilog;
use verilog.vl_types.all;
entity singleCycleProcessor_vlg_vec_tst is
end singleCycleProcessor_vlg_vec_tst;
