    Mac OS X            	   2  �     �                                    ATTR     �    �                    :  com.apple.quarantine   >   H  com.apple.macl FE  �    %com.apple.metadata:kMDItemWhereFroms   �     com.apple.provenance 0281;66101e49;Firefox;DD6BFEED-0585-49F9-A7AF-DA20FF4A9AB1 �B#@AQFO��b^��                                                      bplist00�_khttps://uottawa.brightspace.com/d2l/le/content/417607/topics/files/download/5789974/DirectFileTopicDownload_whttps://uottawa.brightspace.com/d2l/le/content/417607/Home?itemIdentifier=D2L.LE.Content.ContentObject.ModuleCO-5765593y                            �  S���bb                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        This resource fork intentionally left blank                                                                                                                                                                                                                            ��