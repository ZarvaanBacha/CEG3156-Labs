library ieee;
use ieee.std_logic_1164.all;

package utils is
	type matrixnx8 is array(natural range <>) of std_logic_vector(0 to 7);

end package;
