library verilog;
use verilog.vl_types.all;
entity shift_multiplier_8_bit_data_vlg_vec_tst is
end shift_multiplier_8_bit_data_vlg_vec_tst;
