library verilog;
use verilog.vl_types.all;
entity ALUnBit_vlg_vec_tst is
end ALUnBit_vlg_vec_tst;
