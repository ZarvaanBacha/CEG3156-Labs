library verilog;
use verilog.vl_types.all;
entity nBitALU_vlg_vec_tst is
end nBitALU_vlg_vec_tst;
