library verilog;
use verilog.vl_types.all;
entity registerFile_vlg_vec_tst is
end registerFile_vlg_vec_tst;
