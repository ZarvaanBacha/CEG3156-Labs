library verilog;
use verilog.vl_types.all;
entity nBitComparator_vlg_vec_tst is
end nBitComparator_vlg_vec_tst;
