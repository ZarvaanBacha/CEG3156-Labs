library verilog;
use verilog.vl_types.all;
entity DispController_vlg_vec_tst is
end DispController_vlg_vec_tst;
